module furina(input fontaine, input focalor, output celestia);

    assign celestia = fontaine & focalor;

endmodule